// fig_begin hello
module main;

initial
  begin
    $display("Hello, world");
    $finish;
  end

endmodule
// fig_end hello
